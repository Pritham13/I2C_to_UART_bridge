module i2c_tb(); 
reg SCL,SDA; wire [6:0]data;
initial
  begin

endmodule

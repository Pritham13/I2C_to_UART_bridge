module i2c_master(input [7:0]data,
  input clk,
  inout SDA,
  output reg SCL
  );

  always @(posedge clk)
    begin
      
    end
